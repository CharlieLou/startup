module a;
	initial begin
		$display("yeah, this is the beginning\n");
		$display("need color!\n");
	end
endmodule