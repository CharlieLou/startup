module a;
	initial begin
		$display("yeah, this is the beginning\n");
	end
endmodule